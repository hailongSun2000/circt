// RUN:

localparam Z = 9001;
